** sch_path: /home/elastica/resistor_divider_generator/sch/untitled.sch
**.subckt untitled
XR12 net2 net1 net4 sky130_fd_pr__res_xhigh_po_1p41 L=20 mult=1 m=1
XR1 net3 net2 net5 sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR2 net3 net2 net6 sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
**.ends
.end
